----------------------------------------------------------------------------------
-- Company:
-- Engineer:
--
-- Create Date: 15.02.2019 16:46:24
-- Design Name:
-- Module Name: top - Behavioral
-- Project Name:
-- Target Devices:
-- Tool Versions:
-- Description:
--
-- Dependencies:
--
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
----------------------------------------------------------------------------------
LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

ENTITY top IS
	PORT (
		--user pmod
		PMOD_JB : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		PMOD_JC : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		PMOD_JD : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);
		PMOD_JE : INOUT STD_LOGIC_VECTOR(7 DOWNTO 0);

		--clk
		sys_clock : IN STD_LOGIC;
		leds : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);

		--part RGB
		RGB_LED1 : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		RGB_LED2 : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);

		DDR_addr : INOUT STD_LOGIC_VECTOR (14 DOWNTO 0);
		DDR_ba : INOUT STD_LOGIC_VECTOR (2 DOWNTO 0);
		DDR_cas_n : INOUT STD_LOGIC;
		DDR_ck_n : INOUT STD_LOGIC;
		DDR_ck_p : INOUT STD_LOGIC;
		DDR_cke : INOUT STD_LOGIC;
		DDR_cs_n : INOUT STD_LOGIC;
		DDR_dm : INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		DDR_dq : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
		DDR_dqs_n : INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		DDR_dqs_p : INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
		DDR_odt : INOUT STD_LOGIC;
		DDR_ras_n : INOUT STD_LOGIC;
		DDR_reset_n : INOUT STD_LOGIC;
		DDR_we_n : INOUT STD_LOGIC;
		FIXED_IO_ddr_vrn : INOUT STD_LOGIC;
		FIXED_IO_ddr_vrp : INOUT STD_LOGIC;
		FIXED_IO_mio : INOUT STD_LOGIC_VECTOR (53 DOWNTO 0);
		FIXED_IO_ps_clk : INOUT STD_LOGIC;
		FIXED_IO_ps_porb : INOUT STD_LOGIC;
		FIXED_IO_ps_srstb : INOUT STD_LOGIC
	);
END top;

ARCHITECTURE Behavioral OF top IS

    component MUX is
    Port ( 
        SYSCLK_125MHZ : in STD_LOGIC;
        MUX_GPIO : in STD_LOGIC_VECTOR(28 downto 0);
        RGB_LED1 : out STD_LOGIC_VECTOR(2 DOWNTO 0);
        RGB_LED2 : out STD_LOGIC_VECTOR(2 DOWNTO 0);
        LEDS : out STD_LOGIC_VECTOR(3 DOWNTO 0);
               
        PMOD_JB_IN : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OUT : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OE :  out STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JC_IN : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OUT : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OE : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        
        PMOD_JD_IN : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OUT : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OE : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        
        PMOD_JE_IN : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OUT : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OE : out STD_LOGIC_VECTOR(7 DOWNTO 0);
     
        --par0
        PMOD_JB_IN_0 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OUT_0 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OE_0 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JC_IN_0 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OUT_0 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OE_0 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        
        PMOD_JD_IN_0 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OUT_0 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OE_0 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        
        PMOD_JE_IN_0 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OUT_0 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OE_0 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        RGB_LED1_0 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        RGB_LED2_0 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        LEDS_0 : in STD_LOGIC_VECTOR(3 DOWNTO 0);
    
        --par1
        PMOD_JB_IN_1 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OUT_1 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OE_1 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JC_IN_1 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OUT_1 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OE_1 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JD_IN_1 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OUT_1 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OE_1 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JE_IN_1 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OUT_1 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OE_1 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        RGB_LED1_1 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        RGB_LED2_1 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        LEDS_1 : in STD_LOGIC_VECTOR(3 DOWNTO 0);
        --par2
        PMOD_JB_IN_2 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OUT_2 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OE_2 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JC_IN_2 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OUT_2 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OE_2 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JD_IN_2 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OUT_2 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OE_2 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JE_IN_2 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OUT_2 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OE_2 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        RGB_LED1_2 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        RGB_LED2_2 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        LEDS_2 : in STD_LOGIC_VECTOR(3 DOWNTO 0);
    
        --par3
        PMOD_JB_IN_3 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OUT_3 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OE_3 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JC_IN_3 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OUT_3 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OE_3 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JD_IN_3 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OUT_3 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OE_3 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JE_IN_3 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OUT_3 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OE_3 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        RGB_LED1_3 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        RGB_LED2_3 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        LEDS_3 : in STD_LOGIC_VECTOR(3 DOWNTO 0);
    
        --par4
        PMOD_JB_IN_4 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OUT_4 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
         PMOD_JB_OE_4 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JC_IN_4 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OUT_4 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OE_4 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JD_IN_4 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OUT_4 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OE_4 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JE_IN_4 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OUT_4 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OE_4 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        RGB_LED1_4 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        RGB_LED2_4 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        LEDS_4 : in STD_LOGIC_VECTOR(3 DOWNTO 0);
    
        --par5
        PMOD_JB_IN_5 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OUT_5 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OE_5 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JC_IN_5 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OUT_5 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OE_5 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JD_IN_5 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OUT_5 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OE_5 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JE_IN_5 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OUT_5 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OE_5 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        RGB_LED1_5 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        RGB_LED2_5 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        LEDS_5 : in STD_LOGIC_VECTOR(3 DOWNTO 0);
    
        --par6
        PMOD_JB_IN_6 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OUT_6 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OE_6 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JC_IN_6 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OUT_6 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OE_6 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JD_IN_6 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OUT_6 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OE_6 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JE_IN_6 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OUT_6 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OE_6 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        RGB_LED1_6 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        RGB_LED2_6 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        LEDS_6 : in STD_LOGIC_VECTOR(3 DOWNTO 0);
        
        --par7
        PMOD_JB_IN_7 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OUT_7 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JB_OE_7 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JC_IN_7 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OUT_7 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JC_OE_7 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JD_IN_7 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OUT_7 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JD_OE_7 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        PMOD_JE_IN_7 : out STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OUT_7 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
        PMOD_JE_OE_7 : in STD_LOGIC_VECTOR(7 DOWNTO 0);
    
        RGB_LED1_7 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        RGB_LED2_7 : in STD_LOGIC_VECTOR(2 DOWNTO 0);
        LEDS_7 : in STD_LOGIC_VECTOR(3 DOWNTO 0)
       
    );
    end component;


	COMPONENT par0 IS
		PORT (
			CLK_125MHZ : IN STD_LOGIC;
			CLK_MMC : IN STD_LOGIC_VECTOR (0 TO 0);
			CLK_PLL : IN STD_LOGIC_VECTOR (0 TO 0);
 
			reset : IN STD_LOGIC;
 
			PAR_TEST_GPIO0_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO0_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
 
			PMOD_JB_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JC_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JD_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JE_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); 
 
			leds : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
 
			RGB_LED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			RGB_LED2 : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT par1 IS
		PORT (
			CLK_125MHZ : IN STD_LOGIC;
			CLK_MMC : IN STD_LOGIC_VECTOR (0 TO 0);
			CLK_PLL : IN STD_LOGIC_VECTOR (0 TO 0);
 
			reset : IN STD_LOGIC;
 
			PAR_TEST_GPIO0_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO0_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			PMOD_JB_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JC_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JD_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JE_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); 
 
			leds : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
 
			RGB_LED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			RGB_LED2 : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT par2 IS
		PORT (
			CLK_125MHZ : IN STD_LOGIC;
			CLK_MMC : IN STD_LOGIC_VECTOR (0 TO 0);
			CLK_PLL : IN STD_LOGIC_VECTOR (0 TO 0);
 
			reset : IN STD_LOGIC;
 
			PAR_TEST_GPIO0_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO0_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			PMOD_JB_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JC_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JD_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JE_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); 
 
			leds : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
 
			RGB_LED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			RGB_LED2 : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT par3 IS
		PORT (
			CLK_125MHZ : IN STD_LOGIC;
			CLK_MMC : IN STD_LOGIC_VECTOR (0 TO 0);
			CLK_PLL : IN STD_LOGIC_VECTOR (0 TO 0);
 
			reset : IN STD_LOGIC;
 
			PAR_TEST_GPIO0_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO0_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
 
			PMOD_JB_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JC_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JD_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JE_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); 
			leds : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
 
			RGB_LED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			RGB_LED2 : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT par4 IS
		PORT (
			CLK_125MHZ : IN STD_LOGIC;
			CLK_MMC : IN STD_LOGIC_VECTOR (0 TO 0);
			CLK_PLL : IN STD_LOGIC_VECTOR (0 TO 0);
 
			reset : IN STD_LOGIC;
 
			PAR_TEST_GPIO0_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO0_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
 
			PMOD_JB_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JC_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JD_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JE_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); 
			leds : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
 
			RGB_LED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			RGB_LED2 : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT par5 IS
		PORT (
			CLK_125MHZ : IN STD_LOGIC;
			CLK_MMC : IN STD_LOGIC_VECTOR (0 TO 0);
			CLK_PLL : IN STD_LOGIC_VECTOR (0 TO 0);
 
			reset : IN STD_LOGIC;
 
			PAR_TEST_GPIO0_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO0_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
 
			PMOD_JB_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JC_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JD_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JE_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); 
			leds : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
 
			RGB_LED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			RGB_LED2 : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
		);
	END COMPONENT;

	COMPONENT par6 IS
		PORT (
			CLK_125MHZ : IN STD_LOGIC;
			CLK_MMC : IN STD_LOGIC_VECTOR (0 TO 0);
			CLK_PLL : IN STD_LOGIC_VECTOR (0 TO 0);
 
			reset : IN STD_LOGIC;
 
			PAR_TEST_GPIO0_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO0_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
 
			PMOD_JB_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JB_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JC_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JC_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JD_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JD_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
 
			PMOD_JE_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			PMOD_JE_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); 
			leds : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
 
			RGB_LED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			RGB_LED2 : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
		);
	END COMPONENT;
	
	
        COMPONENT par7 IS
            PORT (
                CLK_125MHZ : IN STD_LOGIC;
                CLK_MMC : IN STD_LOGIC_VECTOR (0 TO 0);
                CLK_PLL : IN STD_LOGIC_VECTOR (0 TO 0);
     
                reset : IN STD_LOGIC;
     
                UART_ZYNQ_txd : IN STD_LOGIC;
                UART_ZYNQ_rxd : OUT STD_LOGIC;
     
                PAR_TEST_GPIO0_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
                PAR_TEST_GPIO0_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
     
                PMOD_JB_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
                PMOD_JB_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
                PMOD_JB_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
     
                PMOD_JC_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
                PMOD_JC_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
                PMOD_JC_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
     
                PMOD_JD_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
                PMOD_JD_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
                PMOD_JD_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
     
                PMOD_JE_IN : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
                PMOD_JE_OUT : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
                PMOD_JE_OE : OUT STD_LOGIC_VECTOR(7 DOWNTO 0); 
                leds : OUT STD_LOGIC_VECTOR (3 DOWNTO 0);
     
                RGB_LED : OUT STD_LOGIC_VECTOR (2 DOWNTO 0);
                RGB_LED2 : OUT STD_LOGIC_VECTOR (2 DOWNTO 0)
            );
        END COMPONENT;

	COMPONENT bd_name_wrapper IS
		PORT (
			DDR_cas_n : INOUT STD_LOGIC;
			DDR_cke : INOUT STD_LOGIC;
			DDR_ck_n : INOUT STD_LOGIC;
			DDR_ck_p : INOUT STD_LOGIC;
			DDR_cs_n : INOUT STD_LOGIC;
			DDR_reset_n : INOUT STD_LOGIC;
			DDR_odt : INOUT STD_LOGIC;
			DDR_ras_n : INOUT STD_LOGIC;
			DDR_we_n : INOUT STD_LOGIC;
			DDR_ba : INOUT STD_LOGIC_VECTOR (2 DOWNTO 0);
			DDR_addr : INOUT STD_LOGIC_VECTOR (14 DOWNTO 0);
			DDR_dm : INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			DDR_dq : INOUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			DDR_dqs_n : INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			DDR_dqs_p : INOUT STD_LOGIC_VECTOR (3 DOWNTO 0);
			FIXED_IO_mio : INOUT STD_LOGIC_VECTOR (53 DOWNTO 0);
			FIXED_IO_ddr_vrn : INOUT STD_LOGIC;
			FIXED_IO_ddr_vrp : INOUT STD_LOGIC;
			FIXED_IO_ps_srstb : INOUT STD_LOGIC;
			FIXED_IO_ps_clk : INOUT STD_LOGIC;
			FIXED_IO_ps_porb : INOUT STD_LOGIC;
			UART_ZYNQ_txd : OUT STD_LOGIC;
			UART_ZYNQ_rxd : IN STD_LOGIC;
			CLK_MMC : OUT STD_LOGIC_VECTOR (0 TO 0);
			CLK_PLL : OUT STD_LOGIC_VECTOR (0 TO 0);
			reset_par : OUT STD_LOGIC_VECTOR (15 DOWNTO 0);
			PAR_TEST_GPIO0_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO0_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO1_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO2_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO3_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO4_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO5_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO6_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO7_IN : IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO1_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO2_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO3_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO5_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO6_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO7_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			PAR_TEST_GPIO4_OUT : OUT STD_LOGIC_VECTOR (31 DOWNTO 0);
			MUX_GPO : out STD_LOGIC_VECTOR ( 28 downto 0 )
		);
	END COMPONENT;
 
	COMPONENT OBUF
		PORT (
			I : IN STD_LOGIC;
			O : OUT STD_LOGIC
		);
	END COMPONENT;
 
	COMPONENT IOBUF IS
		PORT (
			I : IN STD_LOGIC;
			O : OUT STD_LOGIC;
			T : IN STD_LOGIC;
			IO : INOUT STD_LOGIC
		);
	END COMPONENT;

	--gpio signals
	SIGNAL reset_par : STD_LOGIC_VECTOR (15 DOWNTO 0);
 
	SIGNAL PAR_TEST_GPIO0_IN_s : STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL PAR_TEST_GPIO0_OUT_s : STD_LOGIC_VECTOR (31 DOWNTO 0);
 
	SIGNAL PAR_TEST_GPIO1_IN : STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL PAR_TEST_GPIO1_OUT : STD_LOGIC_VECTOR (31 DOWNTO 0);
 
	SIGNAL PAR_TEST_GPIO2_IN : STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL PAR_TEST_GPIO2_OUT : STD_LOGIC_VECTOR (31 DOWNTO 0);
 
	SIGNAL PAR_TEST_GPIO3_IN_S : STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL PAR_TEST_GPIO3_OUT_S : STD_LOGIC_VECTOR (31 DOWNTO 0);
 
	SIGNAL PAR_TEST_GPIO4_IN : STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL PAR_TEST_GPIO4_OUT : STD_LOGIC_VECTOR (31 DOWNTO 0);
 
	SIGNAL PAR_TEST_GPIO5_IN : STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL PAR_TEST_GPIO5_OUT : STD_LOGIC_VECTOR (31 DOWNTO 0);
 
	SIGNAL PAR_TEST_GPIO6_IN : STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL PAR_TEST_GPIO6_OUT : STD_LOGIC_VECTOR (31 DOWNTO 0);
 
	SIGNAL PAR_TEST_GPIO7_IN : STD_LOGIC_VECTOR (31 DOWNTO 0);
	SIGNAL PAR_TEST_GPIO7_OUT : STD_LOGIC_VECTOR (31 DOWNTO 0);
 
 
	SIGNAL CLK_MMC : STD_LOGIC_VECTOR(0 DOWNTO 0);
	SIGNAL CLK_PLL : STD_LOGIC_VECTOR(0 DOWNTO 0);
	SIGNAL sys_clk : STD_LOGIC_VECTOR(0 DOWNTO 0);

	SIGNAL UART_ZYNQ_rxd : STD_LOGIC;
	SIGNAL UART_ZYNQ_txd : STD_LOGIC;
 
	SIGNAL PMOD_JB_IN : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OUT : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OE : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JC_IN : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OUT : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OE : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_IN : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OUT : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OE : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_IN : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OUT : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OE : STD_LOGIC_VECTOR(7 DOWNTO 0);
 
	--par0
	SIGNAL PMOD_JB_IN_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OUT_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OE_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JC_IN_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OUT_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OE_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_IN_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OUT_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OE_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_IN_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OUT_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OE_0 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL RGB_LED1_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL RGB_LED2_0 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL LEDS_0 : STD_LOGIC_VECTOR(3 DOWNTO 0);

	--par1
	SIGNAL PMOD_JB_IN_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OUT_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OE_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JC_IN_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OUT_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OE_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JD_IN_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OUT_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OE_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JE_IN_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OUT_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OE_1 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL RGB_LED1_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL RGB_LED2_1 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL LEDS_1 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	--par2
	SIGNAL PMOD_JB_IN_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OUT_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OE_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JC_IN_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OUT_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OE_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JD_IN_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OUT_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OE_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JE_IN_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OUT_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OE_2 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL RGB_LED1_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL RGB_LED2_2 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL LEDS_2 : STD_LOGIC_VECTOR(3 DOWNTO 0);

	--par3
	SIGNAL PMOD_JB_IN_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OUT_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OE_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JC_IN_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OUT_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OE_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JD_IN_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OUT_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OE_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JE_IN_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OUT_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OE_3 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL RGB_LED1_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL RGB_LED2_3 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL LEDS_3 : STD_LOGIC_VECTOR(3 DOWNTO 0);

	--par4
	SIGNAL PMOD_JB_IN_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OUT_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OE_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JC_IN_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OUT_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OE_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JD_IN_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OUT_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OE_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JE_IN_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OUT_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OE_4 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL RGB_LED1_4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL RGB_LED2_4 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL LEDS_4 : STD_LOGIC_VECTOR(3 DOWNTO 0);

	--par5
	SIGNAL PMOD_JB_IN_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OUT_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OE_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JC_IN_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OUT_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OE_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JD_IN_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OUT_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OE_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JE_IN_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OUT_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OE_5 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL RGB_LED1_5 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL RGB_LED2_5 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL LEDS_5 : STD_LOGIC_VECTOR(3 DOWNTO 0);

	--par6
	SIGNAL PMOD_JB_IN_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OUT_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JB_OE_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JC_IN_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OUT_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JC_OE_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JD_IN_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OUT_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JD_OE_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL PMOD_JE_IN_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OUT_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);
	SIGNAL PMOD_JE_OE_6 : STD_LOGIC_VECTOR(7 DOWNTO 0);

	SIGNAL RGB_LED1_6 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL RGB_LED2_6 : STD_LOGIC_VECTOR(2 DOWNTO 0);
	SIGNAL LEDS_6 : STD_LOGIC_VECTOR(3 DOWNTO 0);
	
	--par7
    SIGNAL PMOD_JB_IN_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL PMOD_JB_OUT_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL PMOD_JB_OE_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);

    SIGNAL PMOD_JC_IN_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL PMOD_JC_OUT_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL PMOD_JC_OE_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);

    SIGNAL PMOD_JD_IN_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL PMOD_JD_OUT_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL PMOD_JD_OE_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);

    SIGNAL PMOD_JE_IN_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL PMOD_JE_OUT_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);
    SIGNAL PMOD_JE_OE_7 : STD_LOGIC_VECTOR(7 DOWNTO 0);

    SIGNAL RGB_LED1_7 : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL RGB_LED2_7 : STD_LOGIC_VECTOR(2 DOWNTO 0);
    SIGNAL LEDS_7 : STD_LOGIC_VECTOR(3 DOWNTO 0);

    SIGNAL MUX_GPIO : STD_LOGIC_VECTOR(28 DOWNTO 0);
	SIGNAL RGB_LED_obuf : STD_LOGIC_VECTOR(2 DOWNTO 0);

BEGIN
	bd_name_wrapper_port_map : bd_name_wrapper
	PORT MAP(
		--CLK
		CLK_MMC => CLK_MMC, 
		CLK_PLL => CLK_PLL, 
		 
		--DDR
		DDR_cas_n => DDR_cas_n, 
		DDR_cke => DDR_cke, 
		DDR_ck_n => DDR_ck_n, 
		DDR_ck_p => DDR_ck_p, 
		DDR_cs_n => DDR_cs_n, 
		DDR_reset_n => DDR_reset_n, 
		DDR_odt => DDR_odt, 
		DDR_ras_n => DDR_ras_n, 
		DDR_we_n => DDR_we_n, 
		DDR_ba => DDR_ba, 
		DDR_addr => DDR_addr, 
		DDR_dm => DDR_dm, 
		DDR_dq => DDR_dq, 
		DDR_dqs_n => DDR_dqs_n, 
		DDR_dqs_p => DDR_dqs_p,  
		--FIXEDIO
		FIXED_IO_mio => FIXED_IO_mio, 
		FIXED_IO_ddr_vrn => FIXED_IO_ddr_vrn, 
		FIXED_IO_ddr_vrp => FIXED_IO_ddr_vrp, 
		FIXED_IO_ps_srstb => FIXED_IO_ps_srstb, 
		FIXED_IO_ps_clk => FIXED_IO_ps_clk, 
		FIXED_IO_ps_porb => FIXED_IO_ps_porb, 
 
		--UART
		UART_ZYNQ_txd => UART_ZYNQ_txd, 
		UART_ZYNQ_rxd => UART_ZYNQ_rxd, 
 
		--Shared Reset
		reset_par => reset_par,  
		PAR_TEST_GPIO0_IN => PAR_TEST_GPIO0_IN_s,
		PAR_TEST_GPIO1_IN => PAR_TEST_GPIO1_IN, 
		PAR_TEST_GPIO2_IN => PAR_TEST_GPIO2_IN, 
		PAR_TEST_GPIO3_IN => PAR_TEST_GPIO3_IN_S, 
		PAR_TEST_GPIO4_IN => PAR_TEST_GPIO4_IN, 
		PAR_TEST_GPIO5_IN => PAR_TEST_GPIO5_IN, 
		PAR_TEST_GPIO6_IN => PAR_TEST_GPIO6_IN, 
		PAR_TEST_GPIO7_IN => PAR_TEST_GPIO7_IN, 
 
		PAR_TEST_GPIO0_OUT => PAR_TEST_GPIO0_OUT_s, 
		PAR_TEST_GPIO1_OUT => PAR_TEST_GPIO1_OUT, 
		PAR_TEST_GPIO2_OUT => PAR_TEST_GPIO2_OUT, 
		PAR_TEST_GPIO3_OUT => PAR_TEST_GPIO3_OUT_S, 
		PAR_TEST_GPIO4_OUT => PAR_TEST_GPIO4_OUT,
		PAR_TEST_GPIO5_OUT => PAR_TEST_GPIO5_OUT, 
		PAR_TEST_GPIO6_OUT => PAR_TEST_GPIO6_OUT, 
		PAR_TEST_GPIO7_OUT => PAR_TEST_GPIO7_OUT, 
		
		MUX_GPO => MUX_GPIO
	);
 
	par0pm : par0
	PORT MAP(
		CLK_125MHZ => sys_clock, 
		CLK_MMC => CLK_MMC, 
		CLK_PLL => CLK_PLL, 
 
		reset => reset_par(0), 
 
		PAR_TEST_GPIO0_IN => PAR_TEST_GPIO0_OUT_S, 
		PAR_TEST_GPIO0_OUT => PAR_TEST_GPIO0_IN_S, 
 
		PMOD_JB_IN => PMOD_JB_IN_0, 
		PMOD_JB_OUT => PMOD_JB_OUT_0, 
		PMOD_JB_OE => PMOD_JB_OE_0,
		 
		PMOD_JC_IN => PMOD_JC_IN_0, 
		PMOD_JC_OUT => PMOD_JC_OUT_0, 
		PMOD_JC_OE => PMOD_JC_OE_0, 
 
		PMOD_JD_IN => PMOD_JD_IN_0, 
		PMOD_JD_OUT => PMOD_JD_OUT_0, 
		PMOD_JD_OE => PMOD_JD_OE_0, 
 
		PMOD_JE_IN => PMOD_JE_IN_0, 
		PMOD_JE_OUT => PMOD_JE_OUT_0, 
		PMOD_JE_OE => PMOD_JE_OE_0, 
 
		leds => LEDS_0, 
 
		RGB_LED => RGB_LED1_0, 
		RGB_LED2 => RGB_LED2_0);
 
		par1pm : par1 PORT MAP(
		CLK_125MHZ => sys_clock, 
		CLK_MMC => CLK_MMC, 
		CLK_PLL => CLK_PLL, 
 
		reset => reset_par(1), 
 
		PAR_TEST_GPIO0_IN => PAR_TEST_GPIO1_OUT, 
		PAR_TEST_GPIO0_OUT => PAR_TEST_GPIO1_IN, 
 
		PMOD_JB_IN => PMOD_JB_IN_1, 
		PMOD_JB_OUT => PMOD_JB_OUT_1, 
		PMOD_JB_OE => PMOD_JB_OE_1,
		 
		PMOD_JC_IN => PMOD_JC_IN_1, 
		PMOD_JC_OUT => PMOD_JC_OUT_1, 
		PMOD_JC_OE => PMOD_JC_OE_1, 
 
		PMOD_JD_IN => PMOD_JD_IN_1, 
		PMOD_JD_OUT => PMOD_JD_OUT_1, 
		PMOD_JD_OE => PMOD_JD_OE_1, 
 
		PMOD_JE_IN => PMOD_JE_IN_1, 
		PMOD_JE_OUT => PMOD_JE_OUT_1, 
		PMOD_JE_OE => PMOD_JE_OE_1, 
 
		leds => LEDS_1, 
 
		RGB_LED => RGB_LED1_1, 
		RGB_LED2 => RGB_LED2_1
		);
 
 
		par2pm : par2 PORT MAP(
		CLK_125MHZ => sys_clock, 
		CLK_MMC => CLK_MMC, 
		CLK_PLL => CLK_PLL, 
 
		reset => reset_par(2), 
 
		PAR_TEST_GPIO0_IN => PAR_TEST_GPIO2_OUT, 
		PAR_TEST_GPIO0_OUT => PAR_TEST_GPIO2_IN, 
 
		PMOD_JB_IN => PMOD_JB_IN_2, 
		PMOD_JB_OUT => PMOD_JB_OUT_2, 
		PMOD_JB_OE => PMOD_JB_OE_2,
		 
		PMOD_JC_IN => PMOD_JC_IN_2, 
		PMOD_JC_OUT => PMOD_JC_OUT_2, 
		PMOD_JC_OE => PMOD_JC_OE_2, 
 
		PMOD_JD_IN => PMOD_JD_IN_2, 
		PMOD_JD_OUT => PMOD_JD_OUT_2, 
		PMOD_JD_OE => PMOD_JD_OE_2, 
 
		PMOD_JE_IN => PMOD_JE_IN_2, 
		PMOD_JE_OUT => PMOD_JE_OUT_2, 
		PMOD_JE_OE => PMOD_JE_OE_2, 
 
		leds => LEDS_2, 
 
		RGB_LED => RGB_LED1_2, 
		RGB_LED2 => RGB_LED2_2);
 
		par3pm : par3 PORT MAP(
		CLK_125MHZ => sys_clock, 
		CLK_MMC => CLK_MMC, 
		CLK_PLL => CLK_PLL, 
 
		reset => reset_par(3), 
 
		PAR_TEST_GPIO0_IN => PAR_TEST_GPIO3_OUT_S, 
		PAR_TEST_GPIO0_OUT => PAR_TEST_GPIO3_IN_S, 
 
		PMOD_JB_IN => PMOD_JB_IN_3, 
		PMOD_JB_OUT => PMOD_JB_OUT_3, 
		PMOD_JB_OE => PMOD_JB_OE_3,
		 
		PMOD_JC_IN => PMOD_JC_IN_3, 
		PMOD_JC_OUT => PMOD_JC_OUT_3, 
		PMOD_JC_OE => PMOD_JC_OE_3, 
 
		PMOD_JD_IN => PMOD_JD_IN_3, 
		PMOD_JD_OUT => PMOD_JD_OUT_3, 
		PMOD_JD_OE => PMOD_JD_OE_3, 
 
		PMOD_JE_IN => PMOD_JE_IN_3, 
		PMOD_JE_OUT => PMOD_JE_OUT_3, 
		PMOD_JE_OE => PMOD_JE_OE_3, 
 
		leds => LEDS_3, 
 
		RGB_LED => RGB_LED1_3, 
		RGB_LED2 => RGB_LED2_3);
		
		par4pm : par4 PORT MAP(
		CLK_125MHZ => sys_clock, 
		CLK_MMC => CLK_MMC, 
		CLK_PLL => CLK_PLL, 
 
		reset => reset_par(4), 
 
		PAR_TEST_GPIO0_IN => PAR_TEST_GPIO4_OUT, 
		PAR_TEST_GPIO0_OUT => PAR_TEST_GPIO4_In, 
 
		PMOD_JB_IN => PMOD_JB_IN_4, 
		PMOD_JB_OUT => PMOD_JB_OUT_4, 
		PMOD_JB_OE => PMOD_JB_OE_4,
		 
		PMOD_JC_IN => PMOD_JC_IN_4, 
		PMOD_JC_OUT => PMOD_JC_OUT_4, 
		PMOD_JC_OE => PMOD_JC_OE_4, 
 
		PMOD_JD_IN => PMOD_JD_IN_4, 
		PMOD_JD_OUT => PMOD_JD_OUT_4, 
		PMOD_JD_OE => PMOD_JD_OE_4, 
 
		PMOD_JE_IN => PMOD_JE_IN_4, 
		PMOD_JE_OUT => PMOD_JE_OUT_4, 
		PMOD_JE_OE => PMOD_JE_OE_4, 
 
		leds => LEDS_4, 
 
		RGB_LED => RGB_LED1_4, 
		RGB_LED2 => RGB_LED2_4);
		
		par5pm : par5 PORT MAP(
		CLK_125MHZ => sys_clock, 
		CLK_MMC => CLK_MMC, 
		CLK_PLL => CLK_PLL, 
 
		reset => reset_par(5), 
 
		PAR_TEST_GPIO0_IN => PAR_TEST_GPIO5_OUT, 
		PAR_TEST_GPIO0_OUT => PAR_TEST_GPIO5_IN, 
 
		PMOD_JB_IN => PMOD_JB_IN_5, 
		PMOD_JB_OUT => PMOD_JB_OUT_5, 
		PMOD_JB_OE => PMOD_JB_OE_5
		, 
		PMOD_JC_IN => PMOD_JC_IN_5, 
		PMOD_JC_OUT => PMOD_JC_OUT_5, 
		PMOD_JC_OE => PMOD_JC_OE_5, 
 
		PMOD_JD_IN => PMOD_JD_IN_5, 
		PMOD_JD_OUT => PMOD_JD_OUT_5, 
		PMOD_JD_OE => PMOD_JD_OE_5, 
 
		PMOD_JE_IN => PMOD_JE_IN_5, 
		PMOD_JE_OUT => PMOD_JE_OUT_5, 
		PMOD_JE_OE => PMOD_JE_OE_5, 
 
		leds => LEDS_5, 
 
		RGB_LED => RGB_LED1_5, 
		RGB_LED2 => RGB_LED2_5);

		par6pm : par6 PORT MAP(
		CLK_125MHZ => sys_clock, 
		CLK_MMC => CLK_MMC, 
		CLK_PLL => CLK_PLL, 
  
		reset => reset_par(6), 
 
		PAR_TEST_GPIO0_IN => PAR_TEST_GPIO6_OUT, 
		PAR_TEST_GPIO0_OUT => PAR_TEST_GPIO6_IN, 
 
		PMOD_JB_IN => PMOD_JB_IN_6, 
		PMOD_JB_OUT => PMOD_JB_OUT_6, 
		PMOD_JB_OE => PMOD_JB_OE_6, 
		
		PMOD_JC_IN => PMOD_JC_IN_6, 
		PMOD_JC_OUT => PMOD_JC_OUT_6, 
		PMOD_JC_OE => PMOD_JC_OE_6, 
 
		PMOD_JD_IN => PMOD_JD_IN_6, 
		PMOD_JD_OUT => PMOD_JD_OUT_6, 
		PMOD_JD_OE => PMOD_JD_OE_6, 
 
		PMOD_JE_IN => PMOD_JE_IN_6, 
		PMOD_JE_OUT => PMOD_JE_OUT_6, 
		PMOD_JE_OE => PMOD_JE_OE_6, 
 
		leds => LEDS_6, 
 
		RGB_LED => RGB_LED1_6, 
		RGB_LED2 => RGB_LED2_6);


		par7pm : par7 PORT MAP(
		CLK_125MHZ => sys_clock, 
		CLK_MMC => CLK_MMC, 
		CLK_PLL => CLK_PLL, 
 
		uart_zynq_rxd => uart_zynq_rxd, 
		uart_zynq_txd => uart_zynq_txd, 
		reset => reset_par(7), 
 
		PAR_TEST_GPIO0_IN => PAR_TEST_GPIO7_OUT, 
		PAR_TEST_GPIO0_OUT => PAR_TEST_GPIO7_IN, 
 
		PMOD_JB_IN => PMOD_JB_IN_7, 
		PMOD_JB_OUT => PMOD_JB_OUT_7, 
		PMOD_JB_OE => PMOD_JB_OE_7,
		 
		PMOD_JC_IN => PMOD_JC_IN_7, 
		PMOD_JC_OUT => PMOD_JC_OUT_7, 
		PMOD_JC_OE => PMOD_JC_OE_7, 
 
		PMOD_JD_IN => PMOD_JD_IN_7, 
		PMOD_JD_OUT => PMOD_JD_OUT_7, 
		PMOD_JD_OE => PMOD_JD_OE_7, 
 
		PMOD_JE_IN => PMOD_JE_IN_7, 
		PMOD_JE_OUT => PMOD_JE_OUT_7, 
		PMOD_JE_OE => PMOD_JE_OE_7, 
 
		leds => LEDS_7, 
 
		RGB_LED => RGB_LED1_7, 
		RGB_LED2 => RGB_LED2_7);
		
		
    MUX0: MUX
            Port MAP ( 
                SYSCLK_125MHZ=>sys_clock,
                MUX_GPIO=>MUX_GPIO,
                RGB_LED1=>RGB_LED1,
                RGB_LED2=>RGB_LED2,
                LEDS=>LEDS,
                       
                PMOD_JB_IN=>PMOD_JB_IN,
                PMOD_JB_OUT=>PMOD_JB_OUT,
                PMOD_JB_OE=>PMOD_JB_OE,
            
                PMOD_JC_IN =>PMOD_JC_IN,
                PMOD_JC_OUT=>PMOD_JC_OUT,
                PMOD_JC_OE=>PMOD_JC_OE,
                
                PMOD_JD_IN=>PMOD_JD_IN,
                PMOD_JD_OUT =>PMOD_JD_OUT,
                PMOD_JD_OE=>PMOD_JD_OE,
                
                PMOD_JE_IN=>PMOD_JE_IN,
                PMOD_JE_OUT=>PMOD_JE_OUT,
                PMOD_JE_OE=>PMOD_JE_OE,
             
                --par0
                PMOD_JB_IN_0=>PMOD_JB_IN_0,
                PMOD_JB_OUT_0=>PMOD_JB_OUT_0,
                PMOD_JB_OE_0=>PMOD_JB_OE_0,
            
                PMOD_JC_IN_0=>PMOD_JC_IN_0,
                PMOD_JC_OUT_0=>PMOD_JC_OUT_0,
                PMOD_JC_OE_0=>PMOD_JC_OE_0,
                
                PMOD_JD_IN_0=>PMOD_JD_IN_0,
                PMOD_JD_OUT_0=>PMOD_JD_OUT_0,
                PMOD_JD_OE_0=>PMOD_JD_OE_0,
                
                PMOD_JE_IN_0=>PMOD_JE_IN_0,
                PMOD_JE_OUT_0=>PMOD_JE_OUT_0,
                PMOD_JE_OE_0=>PMOD_JE_OE_0,
            
                RGB_LED1_0=>RGB_LED1_0,
                RGB_LED2_0=>RGB_LED2_0,
                LEDS_0=>LEDS_0,
            
                --par1
                PMOD_JB_IN_1=>PMOD_JB_IN_1,
                PMOD_JB_OUT_1=>PMOD_JB_OUT_1,
                PMOD_JB_OE_1=>PMOD_JB_OE_1,
            
                PMOD_JC_IN_1=>PMOD_JC_IN_1,
                PMOD_JC_OUT_1=>PMOD_JC_OUT_1,
                PMOD_JC_OE_1=>PMOD_JC_OE_1,
            
                PMOD_JD_IN_1=>PMOD_JD_IN_1,
                PMOD_JD_OUT_1=>PMOD_JD_OUT_1,
                PMOD_JD_OE_1=>PMOD_JD_OE_1,
            
                PMOD_JE_IN_1=>PMOD_JE_IN_1,
                PMOD_JE_OUT_1=>PMOD_JE_OUT_1,
                PMOD_JE_OE_1=>PMOD_JE_OE_1,
            
                RGB_LED1_1=>RGB_LED1_1,
                RGB_LED2_1=>RGB_LED2_1,
                LEDS_1=>LEDS_1,
                --par2
                PMOD_JB_IN_2=>PMOD_JB_IN_2,
                PMOD_JB_OUT_2=>PMOD_JB_OUT_2,
                PMOD_JB_OE_2=>PMOD_JB_OE_2,
            
                PMOD_JC_IN_2=>PMOD_JC_IN_2,
                PMOD_JC_OUT_2=>PMOD_JC_OUT_2,
                PMOD_JC_OE_2=>PMOD_JC_OE_2,
            
                PMOD_JD_IN_2=>PMOD_JD_IN_2,
                PMOD_JD_OUT_2=>PMOD_JD_OUT_2,
                PMOD_JD_OE_2=>PMOD_JD_OE_2,
            
                PMOD_JE_IN_2=>PMOD_JE_IN_2,
                PMOD_JE_OUT_2=>PMOD_JE_OUT_2,
                PMOD_JE_OE_2=>PMOD_JE_OE_2,
            
                RGB_LED1_2=>RGB_LED1_2,
                RGB_LED2_2=>RGB_LED2_2,
                LEDS_2=>LEDS_2,
            
                --par3
                PMOD_JB_IN_3=>PMOD_JB_IN_3,
                PMOD_JB_OUT_3=>PMOD_JB_OUT_3,
                PMOD_JB_OE_3=>PMOD_JB_OE_3,
            
                PMOD_JC_IN_3=>PMOD_JC_IN_3,
                PMOD_JC_OUT_3=>PMOD_JC_OUT_3,
                PMOD_JC_OE_3=>PMOD_JC_OE_3,
            
                PMOD_JD_IN_3=>PMOD_JD_IN_3,
                PMOD_JD_OUT_3=>PMOD_JD_OUT_3,
                PMOD_JD_OE_3=>PMOD_JD_OE_3,
            
                PMOD_JE_IN_3=>PMOD_JE_IN_3,
                PMOD_JE_OUT_3=>PMOD_JE_OUT_3,
                PMOD_JE_OE_3=>PMOD_JE_OE_3,
            
                RGB_LED1_3=>RGB_LED1_3,
                RGB_LED2_3=>RGB_LED2_3,
                LEDS_3=>LEDS_3,
            
                --par4
                PMOD_JB_IN_4=>PMOD_JB_IN_4,
                PMOD_JB_OUT_4=>PMOD_JB_OUT_4,
                 PMOD_JB_OE_4=>PMOD_JB_OE_4,
            
                PMOD_JC_IN_4=>PMOD_JC_IN_4,
                PMOD_JC_OUT_4=>PMOD_JC_OUT_4,
                PMOD_JC_OE_4=>PMOD_JC_OE_4,
            
                PMOD_JD_IN_4=>PMOD_JD_IN_4,
                PMOD_JD_OUT_4=>PMOD_JD_OUT_4,
                PMOD_JD_OE_4=>PMOD_JD_OE_4,
            
                PMOD_JE_IN_4=>PMOD_JE_IN_4,
                PMOD_JE_OUT_4=>PMOD_JE_OUT_4,
                PMOD_JE_OE_4=>PMOD_JE_OE_4,
            
                RGB_LED1_4=>RGB_LED1_4,
                RGB_LED2_4=>RGB_LED2_4,
                LEDS_4=>LEDS_4,
            
                --par5
                PMOD_JB_IN_5=>PMOD_JB_IN_5,
                PMOD_JB_OUT_5=>PMOD_JB_OUT_5,
                PMOD_JB_OE_5=>PMOD_JB_OE_5,
            
                PMOD_JC_IN_5=>PMOD_JC_IN_5,
                PMOD_JC_OUT_5=>PMOD_JC_OUT_5,
                PMOD_JC_OE_5=>PMOD_JC_OE_5,
            
                PMOD_JD_IN_5=>PMOD_JD_IN_5,
                PMOD_JD_OUT_5=>PMOD_JD_OUT_5,
                PMOD_JD_OE_5=>PMOD_JD_OE_5,
            
                PMOD_JE_IN_5=>PMOD_JE_IN_5,
                PMOD_JE_OUT_5=>PMOD_JE_OUT_5,
                PMOD_JE_OE_5=>PMOD_JE_OE_5,
            
                RGB_LED1_5=>RGB_LED1_5,
                RGB_LED2_5=>RGB_LED2_5,
                LEDS_5=>LEDS_5,
            
                --par6
                PMOD_JB_IN_6=>PMOD_JB_IN_6,
                PMOD_JB_OUT_6=>PMOD_JB_OUT_6,
                PMOD_JB_OE_6=>PMOD_JB_OE_6,
            
                PMOD_JC_IN_6=>PMOD_JC_IN_6,
                PMOD_JC_OUT_6=>PMOD_JC_OUT_6,
                PMOD_JC_OE_6=>PMOD_JC_OE_6,
            
                PMOD_JD_IN_6=>PMOD_JD_IN_6,
                PMOD_JD_OUT_6=>PMOD_JD_OUT_6,
                PMOD_JD_OE_6=>PMOD_JD_OE_6,
            
                PMOD_JE_IN_6=>PMOD_JE_IN_6,
                PMOD_JE_OUT_6=>PMOD_JE_OUT_6,
                PMOD_JE_OE_6=>PMOD_JE_OE_6,
            
               RGB_LED1_6=>RGB_LED1_6,
                RGB_LED2_6=>RGB_LED2_6,
                LEDS_6=>LEDS_6,
                
                --par7
                PMOD_JB_IN_7=>PMOD_JB_IN_7,
                PMOD_JB_OUT_7=>PMOD_JB_OUT_7,
                PMOD_JB_OE_7=>PMOD_JB_OE_7,
            
                PMOD_JC_IN_7=>PMOD_JC_IN_7,
                PMOD_JC_OUT_7=>PMOD_JC_OUT_7,
                PMOD_JC_OE_7=>PMOD_JC_OE_7,
            
                PMOD_JD_IN_7=>PMOD_JD_IN_7,
                PMOD_JD_OUT_7=>PMOD_JD_OUT_7,
                PMOD_JD_OE_7=>PMOD_JD_OE_7,
            
                PMOD_JE_IN_7=>PMOD_JE_IN_7,
                PMOD_JE_OUT_7=>PMOD_JE_OUT_7,
                PMOD_JE_OE_7=>PMOD_JE_OE_7,
            
                RGB_LED1_7=>RGB_LED1_7,
                RGB_LED2_7=>RGB_LED2_7,
                LEDS_7=>LEDS_7      
            );

	
	IOBUF0 : IOBUF
	PORT MAP(
		I => PMOD_JB_OUT(0), 
		O => PMOD_JB_IN(0), 
		T => PMOD_JB_OE(0), 
		IO => PMOD_JB(0)
	);

	IOBUF1 : IOBUF
	PORT MAP(
		I => PMOD_JB_OUT(1), 
		O => PMOD_JB_IN(1), 
		T => PMOD_JB_OE(1), 
		IO => PMOD_JB(1)
	);

	IOBUF2 : IOBUF
	PORT MAP(
		I => PMOD_JB_OUT(2), 
		O => PMOD_JB_IN(2), 
		T => PMOD_JB_OE(2), 
		IO => PMOD_JB(2)
	);

	IOBUF3 : IOBUF
	PORT MAP(
		I => PMOD_JB_OUT(3), 
		O => PMOD_JB_IN(3), 
		T => PMOD_JB_OE(3), 
		IO => PMOD_JB(3)
	);

	IOBUF4 : IOBUF
	PORT MAP(
		I => PMOD_JB_OUT(4), 
		O => PMOD_JB_IN(4), 
		T => PMOD_JB_OE(4), 
		IO => PMOD_JB(4)
	);

	IOBUF5 : IOBUF
	PORT MAP(
		I => PMOD_JB_OUT(5), 
		O => PMOD_JB_IN(5), 
		T => PMOD_JB_OE(5), 
		IO => PMOD_JB(5)
	);

	IOBUF6 : IOBUF
	PORT MAP(
		I => PMOD_JB_OUT(6), 
		O => PMOD_JB_IN(6), 
		T => PMOD_JB_OE(6), 
		IO => PMOD_JB(6)
	);

	IOBUF7 : IOBUF
	PORT MAP(
		I => PMOD_JB_OUT(7), 
		O => PMOD_JB_IN(7), 
		T => PMOD_JB_OE(7), 
		IO => PMOD_JB(7)
	);
	IOBUF0C : IOBUF
	PORT MAP(
		I => PMOD_JC_OUT(0), 
		O => PMOD_JC_IN(0), 
		T => PMOD_JC_OE(0), 
		IO => PMOD_JC(0)
	);

	IOBUF1C : IOBUF
	PORT MAP(
		I => PMOD_JC_OUT(1), 
		O => PMOD_JC_IN(1), 
		T => PMOD_JC_OE(1), 
		IO => PMOD_JC(1)
	);

	IOBUF2C : IOBUF
	PORT MAP(
		I => PMOD_JC_OUT(2), 
		O => PMOD_JC_IN(2), 
		T => PMOD_JC_OE(2), 
		IO => PMOD_JC(2)
	);

	IOBUF3C : IOBUF
	PORT MAP(
		I => PMOD_JC_OUT(3), 
		O => PMOD_JC_IN(3), 
		T => PMOD_JC_OE(3), 
		IO => PMOD_JC(3)
	);

	IOBUF4C : IOBUF
	PORT MAP(
		I => PMOD_JC_OUT(4), 
		O => PMOD_JC_IN(4), 
		T => PMOD_JC_OE(4), 
		IO => PMOD_JC(4)
	);

	IOBUF5C : IOBUF
	PORT MAP(
		I => PMOD_JC_OUT(5), 
		O => PMOD_JC_IN(5), 
		T => PMOD_JC_OE(5), 
		IO => PMOD_JC(5)
	);

	IOBUF6C : IOBUF
	PORT MAP(
		I => PMOD_JC_OUT(6), 
		O => PMOD_JC_IN(6), 
		T => PMOD_JC_OE(6), 
		IO => PMOD_JC(6)
	);

	IOBUF7C : IOBUF
	PORT MAP(
		I => PMOD_JC_OUT(7), 
		O => PMOD_JC_IN(7), 
		T => PMOD_JC_OE(7), 
		IO => PMOD_JC(7)
	);
	IOBUF0D : IOBUF
	PORT MAP(
		I => PMOD_JD_OUT(0), 
		O => PMOD_JD_IN(0), 
		T => PMOD_JD_OE(0), 
		IO => PMOD_JD(0)
	);

	IOBUF1D : IOBUF
	PORT MAP(
		I => PMOD_JD_OUT(1), 
		O => PMOD_JD_IN(1), 
		T => PMOD_JD_OE(1), 
		IO => PMOD_JD(1)
	);

	IOBUF2D : IOBUF
	PORT MAP(
		I => PMOD_JD_OUT(2), 
		O => PMOD_JD_IN(2), 
		T => PMOD_JD_OE(2), 
		IO => PMOD_JD(2)
	);

	IOBUF3D : IOBUF
	PORT MAP(
		I => PMOD_JD_OUT(3), 
		O => PMOD_JD_IN(3), 
		T => PMOD_JD_OE(3), 
		IO => PMOD_JD(3)
	);

	IOBUF4D : IOBUF
	PORT MAP(
		I => PMOD_JD_OUT(4), 
		O => PMOD_JD_IN(4), 
		T => PMOD_JD_OE(4), 
		IO => PMOD_JD(4)
	);

	IOBUF5D : IOBUF
	PORT MAP(
		I => PMOD_JD_OUT(5), 
		O => PMOD_JD_IN(5), 
		T => PMOD_JD_OE(5), 
		IO => PMOD_JD(5)
	);

	IOBUF6D : IOBUF
	PORT MAP(
		I => PMOD_JD_OUT(6), 
		O => PMOD_JD_IN(6), 
		T => PMOD_JD_OE(6), 
		IO => PMOD_JD(6)
	);

	IOBUF7D : IOBUF
	PORT MAP(
		I => PMOD_JD_OUT(7), 
		O => PMOD_JD_IN(7), 
		T => PMOD_JD_OE(7), 
		IO => PMOD_JD(7)
	);

	IOBUF0E : IOBUF
	PORT MAP(
		I => PMOD_JE_OUT(0), 
		O => PMOD_JE_IN(0), 
		T => PMOD_JE_OE(0), 
		IO => PMOD_JE(0)
	);

	IOBUF1E : IOBUF
	PORT MAP(
		I => PMOD_JE_OUT(1), 
		O => PMOD_JE_IN(1), 
		T => PMOD_JE_OE(1), 
		IO => PMOD_JE(1)
	);

	IOBUF2E : IOBUF
	PORT MAP(
		I => PMOD_JE_OUT(2), 
		O => PMOD_JE_IN(2), 
		T => PMOD_JE_OE(2), 
		IO => PMOD_JE(2)
	);

	IOBUF3E : IOBUF
	PORT MAP(
		I => PMOD_JE_OUT(3), 
		O => PMOD_JE_IN(3), 
		T => PMOD_JE_OE(3), 
		IO => PMOD_JE(3)
	);

	IOBUF4E : IOBUF
	PORT MAP(
		I => PMOD_JE_OUT(4), 
		O => PMOD_JE_IN(4), 
		T => PMOD_JE_OE(4), 
		IO => PMOD_JE(4)
	);

	IOBUF5E : IOBUF
	PORT MAP(
		I => PMOD_JE_OUT(5), 
		O => PMOD_JE_IN(5), 
		T => PMOD_JE_OE(5), 
		IO => PMOD_JE(5)
	);

	IOBUF6E : IOBUF
	PORT MAP(
		I => PMOD_JE_OUT(6), 
		O => PMOD_JE_IN(6), 
		T => PMOD_JE_OE(6), 
		IO => PMOD_JE(6)
	);

	IOBUF7E : IOBUF
	PORT MAP(
		I => PMOD_JE_OUT(7), 
		O => PMOD_JE_IN(7), 
		T => PMOD_JE_OE(7), 
		IO => PMOD_JE(7)
	);

END Behavioral;