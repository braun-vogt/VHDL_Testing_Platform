----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date: 15.02.2019 16:46:24
-- Design Name: 
-- Module Name: top - Behavioral
-- Project Name: 
-- Target Devices: 
-- Tool Versions: 
-- Description: 
-- 
-- Dependencies: 
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
-- 
----------------------------------------------------------------------------------


library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx leaf cells in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity top is
    Port ( CLK : in STD_LOGIC;
           RST : in STD_LOGIC;
           RGB_LED : out STD_LOGIC_VECTOR (2 downto 0));
end top;

architecture Behavioral of top is
component PART is
    Port ( CLK : in STD_LOGIC;
           RST : in STD_LOGIC;
           RGB_LED : out STD_LOGIC_VECTOR (2 downto 0));
end component;
begin
par:part port map(CLK=>clk,rst=>rst,RGB_LED=>RGB_LED);

end Behavioral;
